module sparse_mem();

// your code here


endmodule
