import types_pkg::*;

module sva_container ( 
  input state_values state, 
  input wire[3:0] opcode,
  input clk
  );
                 
//***********************
//  Put assertion code here








endmodule
