`ifndef TEST_COLLECTION__SV
`define TEST_COLLECTION__SV

`include "router_env.sv"

class test_base extends uvm_test;
  `uvm_component_utils(test_base)
  router_env env;

  function new(string name, uvm_component parent);
    super.new(name, parent);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);
    env = router_env::type_id::create("env", this);
  endfunction

//
// The start_of_simulation_phase method from lab1 is moved to final_phase
// for the convinience of seeing the topology and factory registry at the
// end of simulation.  In practice, you should implement both phases to
// display the topology and the factory registry.
//
  virtual function void final_phase(uvm_phase phase);
    super.final_phase(phase);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);
    uvm_top.print_topology();
    factory.print();
  endfunction
endclass

// Lab 2 - Include the packet_da_3.sv file
//
// ToDo
`include "packet_da_3.sv"


class test_da_3_inst extends test_base;
  `uvm_component_utils(test_da_3_inst)

  function new(string name, uvm_component parent);
    super.new(name, parent);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);

    // Lab 2 - Use instance override to configure the packet sequencer
    //         to use packet_da_3 instead of packet
    //
    // ToDo
    set_inst_override_by_type("env.i_agent.seqr.*", packet::get_type(), packet_da_3::get_type());

  endfunction

endclass

// Optional Lab 2 - Create a test to globally set all packet instances to packet_da_3
class test_da_3_type extends test_base;
  `uvm_component_utils(test_da_3_type)
  function new(string name, uvm_component parent);
    super.new(name, parent);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);
    set_type_override_by_type(packet::get_type(), packet_da_3::get_type());
  endfunction
endclass



`endif

