module tb;
    top du();
    initial begin
        #1; 
        $finish;
    end
endmodule