// consumer module here
