module pipe( input [7:0] d_in,
             input clk, valid,
             output reg [7:0] d_out );
reg [7:0] d_1, d_2, d_3;
always @ (posedge clk) begin
  if(valid)
     d_1<= #5 d_in;
  d_2 <= #5 d_1;   
  d_3 <= #5 d_2;   
  d_out<= #5 ~d_3; 
end
endmodule


