library verilog;
use verilog.vl_types.all;
entity test_router is
end test_router;
