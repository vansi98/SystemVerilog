interface router_if(input logic clk);
  import defs::*;
  logic  rst ;
  logic [7:0] valid ;
  logic [7:0] stream ;
  logic [7:0] streamo ;
  logic [7:0] busy ;
  logic [7:0] valido ;
  

endinterface: router_if
