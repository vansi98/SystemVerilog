`ifndef OUTPUT_AGENT__SV
`define OUTPUT_AGENT__SV

// include the oMonitor.sv file
`include "oMonitor.sv"

class output_agent extends uvm_agent;
  // This output agent does not have sequencer and driver, but still require a monitor
  // and the associated port_id,virtual interface and analysis port.
  virtual router_tb_io sigs;          // DUT virtual interface
  int                  port_id = -1;  // Agent's designated port
  oMonitor             mon;
  uvm_analysis_port #(packet) analysis_port;

  `uvm_component_utils_begin(output_agent)
    `uvm_field_int(port_id, UVM_DEFAULT | UVM_DEC)
  `uvm_component_utils_end

  function new(string name, uvm_component parent);
    super.new(name, parent);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);

    mon  = oMonitor::type_id::create("mon", this);

    // The agent retrieves port_id and virtual interface.
    uvm_config_db#(int)::get(this, "", "port_id", port_id);
    uvm_config_db#(virtual router_tb_io)::get(this, "", "sigs", sigs);

    uvm_config_db#(int)::set(this, "*", "port_id", port_id);
    uvm_config_db#(virtual router_tb_io)::set(this, "*", "sigs", sigs);
  endfunction

  virtual function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);

    this.analysis_port = mon.analysis_port;
  endfunction

  virtual function void start_of_simulation_phase(uvm_phase phase);
    super.start_of_simulation_phase(phase);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);
    `uvm_info("AGNTCFG", $sformatf("Using port_id of %0d", port_id), UVM_MEDIUM);
  endfunction: start_of_simulation_phase

endclass

`endif
