// link_if here
