library verilog;
use verilog.vl_types.all;
entity router_if is
    port(
        clock           : in     vl_logic
    );
end router_if;
