`ifndef ROUTER_ENV__SV
`define ROUTER_ENV__SV

`include "input_agent.sv"
`include "reset_agent.sv"

// Lab 4 - Task 9, Step 2
//
// Include the driver_reset_sequence.sv file
//
// ToDo



class router_env extends uvm_env;
  input_agent i_agent;
  reset_agent r_agent;

  `uvm_component_utils(router_env)

  function new(string name, uvm_component parent);
    super.new(name, parent);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    `uvm_info("TRACE", $sformatf("%m"), UVM_HIGH);

    i_agent = input_agent::type_id::create("i_agent", this);
    uvm_config_db #(uvm_object_wrapper)::set(this, "i_agent.seqr.main_phase", "default_sequence", packet_sequence::get_type());
    
    // Lab 4 - Task 9, Step 3
    //
    // Configure i_agent's seqr to execute driver_reset_sequence at reset_phase:
    //
    // uvm_config_db #(uvm_object_wrapper)::set(this, "i_agent.seqr.reset_phase", "default_sequence", driver_reset_sequence::get_type());
    //
    // ToDo



    r_agent = reset_agent::type_id::create("r_agent", this);
    uvm_config_db #(uvm_object_wrapper)::set(this, "r_agent.seqr.reset_phase", "default_sequence", reset_sequence::get_type());

  endfunction

endclass

`endif
