
// create package types here

